module music(clk, addr, data);

// 50 MHz
input clk;
input [12:0] addr;
output [9:0] data;

reg [9:0] data;
reg [9:0] notes [0:1199];

initial begin
	// initialize the notes
	notes[0] =  10'b0000000000;
	notes[1] =  10'b0000000000;
	notes[2] =  10'b0000000000;
	notes[3] =  10'b0000000000;
	notes[4] =  10'b0000000000;
	notes[5] =  10'b0000000000;
	notes[6] =  10'b0000000000;
	notes[7] =  10'b0000000000;
	notes[8] =  10'b0000000000;
	notes[9] =  10'b0000000000;
	notes[10] = 10'b0000000000;
	notes[11] = 10'b0000000000;
	notes[12] = 10'b0000000000;
	notes[13] = 10'b0000000000;
	notes[14] = 10'b0000000000;
	notes[15] = 10'b0000000000;
	notes[16] = 10'b0010000100; // measure 5, start of song
	notes[17] = 10'b0010000100;
	notes[18] = 10'b0000000000;
	notes[19] = 10'b0010000100;
	notes[20] = 10'b0001000010;
	notes[21] = 10'b0000000000;
	notes[22] = 10'b0001000010;
	notes[23] = 10'b0000000000;
	notes[24] = 10'b0100001000; // 6
	notes[25] = 10'b0100001000;
	notes[26] = 10'b0000000000;
	notes[27] = 10'b0100001000;
	notes[28] = 10'b0100001000;
	notes[29] = 10'b0100001000;
	notes[30] = 10'b0000000000;
	notes[31] = 10'b0100001000;
	notes[32] = 10'b0010000100; // 7
	notes[33] = 10'b0010000100;
	notes[34] = 10'b0000000000;
	notes[35] = 10'b0010000100;
	notes[36] = 10'b0001000010;
	notes[37] = 10'b0000000000;
	notes[38] = 10'b0001000010;
	notes[39] = 10'b0000000000;
	notes[40] = 10'b1000010000; // 8
	notes[41] = 10'b1000010000;
	notes[42] = 10'b0000000000;
	notes[43] = 10'b1000010000;
	notes[44] = 10'b1000010000;
	notes[45] = 10'b1000010000;
	notes[46] = 10'b0000000000;
	notes[47] = 10'b0000000000;
	notes[48] = 10'b0010000100; // 9
	notes[49] = 10'b0010000100;
	notes[50] = 10'b0000000000;
	notes[51] = 10'b0010000100;
	notes[52] = 10'b0001000010;
	notes[53] = 10'b0000000000;
	notes[54] = 10'b0001000010;
	notes[55] = 10'b0000000000;
	notes[56] = 10'b0100001000; // 10
	notes[57] = 10'b0100001000;
	notes[58] = 10'b0000000000;
	notes[59] = 10'b0100001000;
	notes[60] = 10'b0100001000;
	notes[61] = 10'b0100001000;
	notes[62] = 10'b0000000000;
	notes[63] = 10'b0100001000;
	notes[64] = 10'b0010000100; // 11
	notes[65] = 10'b0010000100;
	notes[66] = 10'b0000000000;
	notes[67] = 10'b0010000100;
	notes[68] = 10'b0001000010;
	notes[69] = 10'b0000000000;
	notes[70] = 10'b0001000010;
	notes[71] = 10'b0000000000;
	notes[72] = 10'b0010010000; // 12
	notes[73] = 10'b0010001000;
	notes[74] = 10'b0010000100;
	notes[75] = 10'b0010000000;
	notes[76] = 10'b0100000100;
	notes[77] = 10'b0100000010;
	notes[78] = 10'b0100000010;
	notes[79] = 10'b0100000000;
	notes[80] = 10'b0010001100; // 13
	notes[81] = 10'b0010001100;
	notes[82] = 10'b0000000000;
	notes[83] = 10'b0010000100;
	notes[84] = 10'b0001000010;
	notes[85] = 10'b0000000000;
	notes[86] = 10'b0001000010;
	notes[87] = 10'b0000000000;
	notes[88] = 10'b0100010100; // 14
	notes[89] = 10'b0100010100;
	notes[90] = 10'b0000000000;
	notes[91] = 10'b0100010100;
	notes[92] = 10'b0100010100;
	notes[93] = 10'b0100010100;
	notes[94] = 10'b0000000000;
	notes[95] = 10'b0100010100;
	notes[96] = 10'b0010001100; // 15
	notes[97] = 10'b0010001100;
	notes[98] = 10'b0000000000;
	notes[99] = 10'b0010000100;
	notes[100] = 10'b0001000010;
	notes[101] = 10'b0000000000;
	notes[102] = 10'b0001000010;
	notes[103] = 10'b0000000000;
	notes[104] = 10'b1000011000; // 16
	notes[105] = 10'b1000011000;
	notes[106] = 10'b0000000000;
	notes[107] = 10'b1000011000;
	notes[108] = 10'b1000011000;
	notes[109] = 10'b1000011000;
	notes[110] = 10'b0000000000;
	notes[111] = 10'b0000011000;
	notes[112] = 10'b0010001100; // 17
	notes[113] = 10'b0010001100;
	notes[114] = 10'b0000000000;
	notes[115] = 10'b0010000100;
	notes[116] = 10'b0001000010;
	notes[117] = 10'b0000000000;
	notes[118] = 10'b0001000010;
	notes[119] = 10'b0000000000;
	notes[120] = 10'b0100010100; // 18
	notes[121] = 10'b0100010100;
	notes[122] = 10'b0000000000;
	notes[123] = 10'b0100010100;
	notes[124] = 10'b0100010100;
	notes[125] = 10'b0100010100;
	notes[126] = 10'b0000000000;
	notes[127] = 10'b0100010100;
	notes[128] = 10'b0010001100; // 19
	notes[129] = 10'b0010001100;
	notes[130] = 10'b0000000000;
	notes[131] = 10'b0010000100;
	notes[132] = 10'b0001000010;
	notes[133] = 10'b0000000000;
	notes[134] = 10'b0001000010;
	notes[135] = 10'b0000000000;
	notes[136] = 10'b0010001010; // 20
	notes[137] = 10'b0010001010;
	notes[138] = 10'b0010001010;
	notes[139] = 10'b0010000000;
	notes[140] = 10'b0100001100;
	notes[141] = 10'b0100001100;
	notes[142] = 10'b0100001100;
	notes[143] = 10'b0000000000;
	notes[144] = 10'b0010001000; // 21
	notes[145] = 10'b0010000000;
	notes[146] = 10'b0000001000;
	notes[147] = 10'b0010001000;
	notes[148] = 10'b0001001000;
	notes[149] = 10'b0000000100;
	notes[150] = 10'b0001001000;
	notes[151] = 10'b0000000100;
	notes[152] = 10'b0100001000; // 22
	notes[153] = 10'b0100000000;
	notes[154] = 10'b0000001000;
	notes[155] = 10'b0100001000;
	notes[156] = 10'b0100001000;
	notes[157] = 10'b0100000100;
	notes[158] = 10'b0000001000;
	notes[159] = 10'b0100000100;
	notes[160] = 10'b0010001000; // 23
	notes[161] = 10'b0010000000;
	notes[162] = 10'b0000001000;
	notes[163] = 10'b0010001000;
	notes[164] = 10'b0001001000;
	notes[165] = 10'b0000000100;
	notes[166] = 10'b0001001000;
	notes[167] = 10'b0000000100;
	notes[168] = 10'b1000001000; // 24
	notes[169] = 10'b1000000000;
	notes[170] = 10'b0000001000;
	notes[171] = 10'b1000001000;
	notes[172] = 10'b1000001000;
	notes[173] = 10'b1000010000;
	notes[174] = 10'b0000010000;
	notes[175] = 10'b0000010000;
	notes[176] = 10'b0010001000; // 25
	notes[177] = 10'b0010000000;
	notes[178] = 10'b0000001000;
	notes[179] = 10'b0010001000;
	notes[180] = 10'b0001001000;
	notes[181] = 10'b0000000100;
	notes[182] = 10'b0001001000;
	notes[183] = 10'b0000000100;
	notes[184] = 10'b0100001000; // 26
	notes[185] = 10'b0100000000;
	notes[1199] = 10'b0000000000;

end

always @(posedge clk) begin
	// give data
	data = notes[addr];
end
endmodule

